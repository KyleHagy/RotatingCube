module RotationOfCube(PointsDrawLine, 
                        VertexBuffer,
                        RotatedVertexBuffer, 
                        FrameBuffer,
                        );

  parameter ROTATE_AXIS = 0;
  parameter THETA = 0;
  parameter SIZE = 0;
  parameter VERTEX_POINT = 0;

  output logic [15:0] PointsDrawLine[11:0][1:0];
  output logic signed [15:0] VertexBuffer[8][3];
  output logic signed [15:0] RotatedVertexBuffer[8][3];
  output logic FrameBuffer[SIZE:0][SIZE:0];


  localparam ROTATE_Z = 0;
  localparam ROTATE_Y = 1;
  localparam ROTATE_X = 2;
  localparam ROTATE_ALL = 3;


  reg signed [31:0] sin[180:0];
  reg signed [31:0] cos[180:0]; 

  reg signed [31:0]sinTheta;  //EX: 32'b0000000000000000_1011010100000100;
  reg signed [31:0]cosTheta;

  reg signed [31:0] cordX;
  reg signed [31:0] cordY;  
  reg signed [31:0] cordZ;   

  reg signed [63:0] XsinTheta;
  reg signed [63:0] XcosTheta;
  reg signed [63:0] YsinTheta;
  reg signed [63:0] YcosTheta;
  reg signed [63:0] ZsinTheta;
  reg signed [63:0] ZcosTheta;

  integer newCordX;
  integer newCordY;
  integer newCordZ;



  integer x1, x2, y1, y2, z1, z2;
  integer xs, dx, dxAbs;
  integer ys, dy, dyAbs;
  integer zs, dz, dzAbs;
  integer p1, p2;
  

  always @(*) begin
    
    sin[0] = 32'b0000000000000000_0000000000000000;
    sin[1] = 32'b0000000000000000_0000010001110111;
    sin[2] = 32'b0000000000000000_0000100011101111;
    sin[3] = 32'b0000000000000000_0000110101100101;
    sin[4] = 32'b0000000000000000_0001000111011011;
    sin[5] = 32'b0000000000000000_0001011001001111;
    sin[6] = 32'b0000000000000000_0001101011000010;
    sin[7] = 32'b0000000000000000_0001111100110010;
    sin[8] = 32'b0000000000000000_0010001110100000;
    sin[9] = 32'b0000000000000000_0010100000001100;
    sin[10] = 32'b0000000000000000_0010110001110100;
    sin[11] = 32'b0000000000000000_0011000011011000;
    sin[12] = 32'b0000000000000000_0011010100111001;
    sin[13] = 32'b0000000000000000_0011100110010110;
    sin[14] = 32'b0000000000000000_0011110111101110;
    sin[15] = 32'b0000000000000000_0100001001000001;
    sin[16] = 32'b0000000000000000_0100011010010000;
    sin[17] = 32'b0000000000000000_0100101011011000;
    sin[18] = 32'b0000000000000000_0100111100011011;
    sin[19] = 32'b0000000000000000_0101001101011000;
    sin[20] = 32'b0000000000000000_0101011110001110;
    sin[21] = 32'b0000000000000000_0101101110111110;
    sin[22] = 32'b0000000000000000_0101111111100110;
    sin[23] = 32'b0000000000000000_0110010000000110;
    sin[24] = 32'b0000000000000000_0110100000011111;
    sin[25] = 32'b0000000000000000_0110110000110000;
    sin[26] = 32'b0000000000000000_0111000000111001;
    sin[27] = 32'b0000000000000000_0111010000111000;
    sin[28] = 32'b0000000000000000_0111100000101111;
    sin[29] = 32'b0000000000000000_0111110000011100;
    sin[30] = 32'b0000000000000000_0111111111111111;
    sin[31] = 32'b0000000000000000_1000001111011001;
    sin[32] = 32'b0000000000000000_1000011110101000;
    sin[33] = 32'b0000000000000000_1000101101101101;
    sin[34] = 32'b0000000000000000_1000111100100111;
    sin[35] = 32'b0000000000000000_1001001011010101;
    sin[36] = 32'b0000000000000000_1001011001111001;
    sin[37] = 32'b0000000000000000_1001101000010000;
    sin[38] = 32'b0000000000000000_1001110110011011;
    sin[39] = 32'b0000000000000000_1010000100011011;
    sin[40] = 32'b0000000000000000_1010010010001101;
    sin[41] = 32'b0000000000000000_1010011111110011;
    sin[42] = 32'b0000000000000000_1010101101001100;
    sin[43] = 32'b0000000000000000_1010111010010111;
    sin[44] = 32'b0000000000000000_1011000111010101;
    sin[45] = 32'b0000000000000000_1011010100000100;
    sin[46] = 32'b0000000000000000_1011100000100110;
    sin[47] = 32'b0000000000000000_1011101100111001;
    sin[48] = 32'b0000000000000000_1011111000111110;
    sin[49] = 32'b0000000000000000_1100000100110100;
    sin[50] = 32'b0000000000000000_1100010000011011;
    sin[51] = 32'b0000000000000000_1100011011110011;
    sin[52] = 32'b0000000000000000_1100100110111011;
    sin[53] = 32'b0000000000000000_1100110001110011;
    sin[54] = 32'b0000000000000000_1100111100011011;
    sin[55] = 32'b0000000000000000_1101000110110011;
    sin[56] = 32'b0000000000000000_1101010000111011;
    sin[57] = 32'b0000000000000000_1101011010110011;
    sin[58] = 32'b0000000000000000_1101100100011001;
    sin[59] = 32'b0000000000000000_1101101101101111;
    sin[60] = 32'b0000000000000000_1101110110110011;
    sin[61] = 32'b0000000000000000_1101111111100111;
    sin[62] = 32'b0000000000000000_1110001000001000;
    sin[63] = 32'b0000000000000000_1110010000011001;
    sin[64] = 32'b0000000000000000_1110011000010111;
    sin[65] = 32'b0000000000000000_1110100000000011;
    sin[66] = 32'b0000000000000000_1110100111011110;
    sin[67] = 32'b0000000000000000_1110101110100110;
    sin[68] = 32'b0000000000000000_1110110101011011;
    sin[69] = 32'b0000000000000000_1110111011111111;
    sin[70] = 32'b0000000000000000_1111000010001111;
    sin[71] = 32'b0000000000000000_1111001000001101;
    sin[72] = 32'b0000000000000000_1111001101111000;
    sin[73] = 32'b0000000000000000_1111010011010000;
    sin[74] = 32'b0000000000000000_1111011000010101;
    sin[75] = 32'b0000000000000000_1111011101000110;
    sin[76] = 32'b0000000000000000_1111100001100101;
    sin[77] = 32'b0000000000000000_1111100101110000;
    sin[78] = 32'b0000000000000000_1111101001100111;
    sin[79] = 32'b0000000000000000_1111101101001011;
    sin[80] = 32'b0000000000000000_1111110000011100;
    sin[81] = 32'b0000000000000000_1111110011011001;
    sin[82] = 32'b0000000000000000_1111110110000010;
    sin[83] = 32'b0000000000000000_1111111000010111;
    sin[84] = 32'b0000000000000000_1111111010011000;
    sin[85] = 32'b0000000000000000_1111111100000110;
    sin[86] = 32'b0000000000000000_1111111101100000;
    sin[87] = 32'b0000000000000000_1111111110100110;
    sin[88] = 32'b0000000000000000_1111111111011000;
    sin[89] = 32'b0000000000000000_1111111111110110;
    sin[90] = 32'b0000000000000001_0000000000000000;
    sin[91] = 32'b0000000000000000_1111111111110110;
    sin[92] = 32'b0000000000000000_1111111111011000;
    sin[93] = 32'b0000000000000000_1111111110100110;
    sin[94] = 32'b0000000000000000_1111111101100000;
    sin[95] = 32'b0000000000000000_1111111100000110;
    sin[96] = 32'b0000000000000000_1111111010011000;
    sin[97] = 32'b0000000000000000_1111111000010111;
    sin[98] = 32'b0000000000000000_1111110110000010;
    sin[99] = 32'b0000000000000000_1111110011011001;
    sin[100] = 32'b0000000000000000_1111110000011100;
    sin[101] = 32'b0000000000000000_1111101101001011;
    sin[102] = 32'b0000000000000000_1111101001100111;
    sin[103] = 32'b0000000000000000_1111100101110000;
    sin[104] = 32'b0000000000000000_1111100001100101;
    sin[105] = 32'b0000000000000000_1111011101000110;
    sin[106] = 32'b0000000000000000_1111011000010101;
    sin[107] = 32'b0000000000000000_1111010011010000;
    sin[108] = 32'b0000000000000000_1111001101111000;
    sin[109] = 32'b0000000000000000_1111001000001101;
    sin[110] = 32'b0000000000000000_1111000010001111;
    sin[111] = 32'b0000000000000000_1110111011111111;
    sin[112] = 32'b0000000000000000_1110110101011011;
    sin[113] = 32'b0000000000000000_1110101110100110;
    sin[114] = 32'b0000000000000000_1110100111011110;
    sin[115] = 32'b0000000000000000_1110100000000011;
    sin[116] = 32'b0000000000000000_1110011000010111;
    sin[117] = 32'b0000000000000000_1110010000011001;
    sin[118] = 32'b0000000000000000_1110001000001000;
    sin[119] = 32'b0000000000000000_1101111111100111;
    sin[120] = 32'b0000000000000000_1101110110110011;
    sin[121] = 32'b0000000000000000_1101101101101111;
    sin[122] = 32'b0000000000000000_1101100100011001;
    sin[123] = 32'b0000000000000000_1101011010110011;
    sin[124] = 32'b0000000000000000_1101010000111011;
    sin[125] = 32'b0000000000000000_1101000110110011;
    sin[126] = 32'b0000000000000000_1100111100011011;
    sin[127] = 32'b0000000000000000_1100110001110011;
    sin[128] = 32'b0000000000000000_1100100110111011;
    sin[129] = 32'b0000000000000000_1100011011110011;
    sin[130] = 32'b0000000000000000_1100010000011011;
    sin[131] = 32'b0000000000000000_1100000100110100;
    sin[132] = 32'b0000000000000000_1011111000111110;
    sin[133] = 32'b0000000000000000_1011101100111001;
    sin[134] = 32'b0000000000000000_1011100000100110;
    sin[135] = 32'b0000000000000000_1011010100000100;
    sin[136] = 32'b0000000000000000_1011000111010101;
    sin[137] = 32'b0000000000000000_1010111010010111;
    sin[138] = 32'b0000000000000000_1010101101001100;
    sin[139] = 32'b0000000000000000_1010011111110011;
    sin[140] = 32'b0000000000000000_1010010010001101;
    sin[141] = 32'b0000000000000000_1010000100011011;
    sin[142] = 32'b0000000000000000_1001110110011011;
    sin[143] = 32'b0000000000000000_1001101000010000;
    sin[144] = 32'b0000000000000000_1001011001111001;
    sin[145] = 32'b0000000000000000_1001001011010101;
    sin[146] = 32'b0000000000000000_1000111100100111;
    sin[147] = 32'b0000000000000000_1000101101101101;
    sin[148] = 32'b0000000000000000_1000011110101000;
    sin[149] = 32'b0000000000000000_1000001111011001;
    sin[150] = 32'b0000000000000000_0111111111111111;
    sin[151] = 32'b0000000000000000_0111110000011100;
    sin[152] = 32'b0000000000000000_0111100000101111;
    sin[153] = 32'b0000000000000000_0111010000111000;
    sin[154] = 32'b0000000000000000_0111000000111001;
    sin[155] = 32'b0000000000000000_0110110000110000;
    sin[156] = 32'b0000000000000000_0110100000011111;
    sin[157] = 32'b0000000000000000_0110010000000110;
    sin[158] = 32'b0000000000000000_0101111111100110;
    sin[159] = 32'b0000000000000000_0101101110111110;
    sin[160] = 32'b0000000000000000_0101011110001110;
    sin[161] = 32'b0000000000000000_0101001101011000;
    sin[162] = 32'b0000000000000000_0100111100011011;
    sin[163] = 32'b0000000000000000_0100101011011000;
    sin[164] = 32'b0000000000000000_0100011010010000;
    sin[165] = 32'b0000000000000000_0100001001000001;
    sin[166] = 32'b0000000000000000_0011110111101110;
    sin[167] = 32'b0000000000000000_0011100110010110;
    sin[168] = 32'b0000000000000000_0011010100111001;
    sin[169] = 32'b0000000000000000_0011000011011000;
    sin[170] = 32'b0000000000000000_0010110001110100;
    sin[171] = 32'b0000000000000000_0010100000001100;
    sin[172] = 32'b0000000000000000_0010001110100000;
    sin[173] = 32'b0000000000000000_0001111100110010;
    sin[174] = 32'b0000000000000000_0001101011000010;
    sin[175] = 32'b0000000000000000_0001011001001111;
    sin[176] = 32'b0000000000000000_0001000111011011;
    sin[177] = 32'b0000000000000000_0000110101100101;
    sin[178] = 32'b0000000000000000_0000100011101111;
    sin[179] = 32'b0000000000000000_0000010001110111;
    sin[180] = 32'b0000000000000000_0000000000000000;




    cos[0] = 32'b0000000000000001_0000000000000000;
    cos[1] = 32'b0000000000000000_1111111111110110;
    cos[2] = 32'b0000000000000000_1111111111011000;
    cos[3] = 32'b0000000000000000_1111111110100110;
    cos[4] = 32'b0000000000000000_1111111101100000;
    cos[5] = 32'b0000000000000000_1111111100000110;
    cos[6] = 32'b0000000000000000_1111111010011000;
    cos[7] = 32'b0000000000000000_1111111000010111;
    cos[8] = 32'b0000000000000000_1111110110000010;
    cos[9] = 32'b0000000000000000_1111110011011001;
    cos[10] = 32'b0000000000000000_1111110000011100;
    cos[11] = 32'b0000000000000000_1111101101001011;
    cos[12] = 32'b0000000000000000_1111101001100111;
    cos[13] = 32'b0000000000000000_1111100101110000;
    cos[14] = 32'b0000000000000000_1111100001100101;
    cos[15] = 32'b0000000000000000_1111011101000110;
    cos[16] = 32'b0000000000000000_1111011000010101;
    cos[17] = 32'b0000000000000000_1111010011010000;
    cos[18] = 32'b0000000000000000_1111001101111000;
    cos[19] = 32'b0000000000000000_1111001000001101;
    cos[20] = 32'b0000000000000000_1111000010001111;
    cos[21] = 32'b0000000000000000_1110111011111111;
    cos[22] = 32'b0000000000000000_1110110101011011;
    cos[23] = 32'b0000000000000000_1110101110100110;
    cos[24] = 32'b0000000000000000_1110100111011110;
    cos[25] = 32'b0000000000000000_1110100000000011;
    cos[26] = 32'b0000000000000000_1110011000010111;
    cos[27] = 32'b0000000000000000_1110010000011001;
    cos[28] = 32'b0000000000000000_1110001000001000;
    cos[29] = 32'b0000000000000000_1101111111100111;
    cos[30] = 32'b0000000000000000_1101110110110011;
    cos[31] = 32'b0000000000000000_1101101101101111;
    cos[32] = 32'b0000000000000000_1101100100011001;
    cos[33] = 32'b0000000000000000_1101011010110011;
    cos[34] = 32'b0000000000000000_1101010000111011;
    cos[35] = 32'b0000000000000000_1101000110110011;
    cos[36] = 32'b0000000000000000_1100111100011011;
    cos[37] = 32'b0000000000000000_1100110001110011;
    cos[38] = 32'b0000000000000000_1100100110111011;
    cos[39] = 32'b0000000000000000_1100011011110011;
    cos[40] = 32'b0000000000000000_1100010000011011;
    cos[41] = 32'b0000000000000000_1100000100110100;
    cos[42] = 32'b0000000000000000_1011111000111110;
    cos[43] = 32'b0000000000000000_1011101100111001;
    cos[44] = 32'b0000000000000000_1011100000100110;
    cos[45] = 32'b0000000000000000_1011010100000100;
    cos[46] = 32'b0000000000000000_1011000111010101;
    cos[47] = 32'b0000000000000000_1010111010010111;
    cos[48] = 32'b0000000000000000_1010101101001100;
    cos[49] = 32'b0000000000000000_1010011111110011;
    cos[50] = 32'b0000000000000000_1010010010001101;
    cos[51] = 32'b0000000000000000_1010000100011011;
    cos[52] = 32'b0000000000000000_1001110110011011;
    cos[53] = 32'b0000000000000000_1001101000010000;
    cos[54] = 32'b0000000000000000_1001011001111001;
    cos[55] = 32'b0000000000000000_1001001011010101;
    cos[56] = 32'b0000000000000000_1000111100100111;
    cos[57] = 32'b0000000000000000_1000101101101101;
    cos[58] = 32'b0000000000000000_1000011110101000;
    cos[59] = 32'b0000000000000000_1000001111011001;
    cos[60] = 32'b0000000000000000_1000000000000000;
    cos[61] = 32'b0000000000000000_0111110000011100;
    cos[62] = 32'b0000000000000000_0111100000101111;
    cos[63] = 32'b0000000000000000_0111010000111000;
    cos[64] = 32'b0000000000000000_0111000000111001;
    cos[65] = 32'b0000000000000000_0110110000110000;
    cos[66] = 32'b0000000000000000_0110100000011111;
    cos[67] = 32'b0000000000000000_0110010000000110;
    cos[68] = 32'b0000000000000000_0101111111100110;
    cos[69] = 32'b0000000000000000_0101101110111110;
    cos[70] = 32'b0000000000000000_0101011110001110;
    cos[71] = 32'b0000000000000000_0101001101011000;
    cos[72] = 32'b0000000000000000_0100111100011011;
    cos[73] = 32'b0000000000000000_0100101011011000;
    cos[74] = 32'b0000000000000000_0100011010010000;
    cos[75] = 32'b0000000000000000_0100001001000001;
    cos[76] = 32'b0000000000000000_0011110111101110;
    cos[77] = 32'b0000000000000000_0011100110010110;
    cos[78] = 32'b0000000000000000_0011010100111001;
    cos[79] = 32'b0000000000000000_0011000011011000;
    cos[80] = 32'b0000000000000000_0010110001110100;
    cos[81] = 32'b0000000000000000_0010100000001100;
    cos[82] = 32'b0000000000000000_0010001110100000;
    cos[83] = 32'b0000000000000000_0001111100110010;
    cos[84] = 32'b0000000000000000_0001101011000010;
    cos[85] = 32'b0000000000000000_0001011001001111;
    cos[86] = 32'b0000000000000000_0001000111011011;
    cos[87] = 32'b0000000000000000_0000110101100101;
    cos[88] = 32'b0000000000000000_0000100011101111;
    cos[89] = 32'b0000000000000000_0000010001110111;
    cos[90] = 32'b0000000000000000_0000000000000000;
    cos[91] = 32'b1111111111111111_1111101110001001;
    cos[92] = 32'b1111111111111111_1111011100010001;
    cos[93] = 32'b1111111111111111_1111001010011011;
    cos[94] = 32'b1111111111111111_1110111000100101;
    cos[95] = 32'b1111111111111111_1110100110110001;
    cos[96] = 32'b1111111111111111_1110010100111110;
    cos[97] = 32'b1111111111111111_1110000011001110;
    cos[98] = 32'b1111111111111111_1101110001100000;
    cos[99] = 32'b1111111111111111_1101011111110100;
    cos[100] = 32'b1111111111111111_1101001110001100;
    cos[101] = 32'b1111111111111111_1100111100101000;
    cos[102] = 32'b1111111111111111_1100101011000111;
    cos[103] = 32'b1111111111111111_1100011001101010;
    cos[104] = 32'b1111111111111111_1100001000010010;
    cos[105] = 32'b1111111111111111_1011110110111111;
    cos[106] = 32'b1111111111111111_1011100101110000;
    cos[107] = 32'b1111111111111111_1011010100101000;
    cos[108] = 32'b1111111111111111_1011000011100101;
    cos[109] = 32'b1111111111111111_1010110010101000;
    cos[110] = 32'b1111111111111111_1010100001110010;
    cos[111] = 32'b1111111111111111_1010010001000010;
    cos[112] = 32'b1111111111111111_1010000000011010;
    cos[113] = 32'b1111111111111111_1001101111111010;
    cos[114] = 32'b1111111111111111_1001011111100001;
    cos[115] = 32'b1111111111111111_1001001111010000;
    cos[116] = 32'b1111111111111111_1000111111000111;
    cos[117] = 32'b1111111111111111_1000101111001000;
    cos[118] = 32'b1111111111111111_1000011111010001;
    cos[119] = 32'b1111111111111111_1000001111100100;
    cos[120] = 32'b1111111111111111_1000000000000000;
    cos[121] = 32'b1111111111111111_0111110000100111;
    cos[122] = 32'b1111111111111111_0111100001011000;
    cos[123] = 32'b1111111111111111_0111010010010011;
    cos[124] = 32'b1111111111111111_0111000011011001;
    cos[125] = 32'b1111111111111111_0110110100101011;
    cos[126] = 32'b1111111111111111_0110100110000111;
    cos[127] = 32'b1111111111111111_0110010111110000;
    cos[128] = 32'b1111111111111111_0110001001100101;
    cos[129] = 32'b1111111111111111_0101111011100101;
    cos[130] = 32'b1111111111111111_0101101101110011;
    cos[131] = 32'b1111111111111111_0101100000001101;
    cos[132] = 32'b1111111111111111_0101010010110100;
    cos[133] = 32'b1111111111111111_0101000101101001;
    cos[134] = 32'b1111111111111111_0100111000101011;
    cos[135] = 32'b1111111111111111_0100101011111100;
    cos[136] = 32'b1111111111111111_0100011111011010;
    cos[137] = 32'b1111111111111111_0100010011000111;
    cos[138] = 32'b1111111111111111_0100000111000010;
    cos[139] = 32'b1111111111111111_0011111011001100;
    cos[140] = 32'b1111111111111111_0011101111100101;
    cos[141] = 32'b1111111111111111_0011100100001101;
    cos[142] = 32'b1111111111111111_0011011001000101;
    cos[143] = 32'b1111111111111111_0011001110001101;
    cos[144] = 32'b1111111111111111_0011000011100101;
    cos[145] = 32'b1111111111111111_0010111001001101;
    cos[146] = 32'b1111111111111111_0010101111000101;
    cos[147] = 32'b1111111111111111_0010100101001101;
    cos[148] = 32'b1111111111111111_0010011011100111;
    cos[149] = 32'b1111111111111111_0010010010010001;
    cos[150] = 32'b1111111111111111_0010001001001101;
    cos[151] = 32'b1111111111111111_0010000000011001;
    cos[152] = 32'b1111111111111111_0001110111111000;
    cos[153] = 32'b1111111111111111_0001101111100111;
    cos[154] = 32'b1111111111111111_0001100111101001;
    cos[155] = 32'b1111111111111111_0001011111111101;
    cos[156] = 32'b1111111111111111_0001011000100010;
    cos[157] = 32'b1111111111111111_0001010001011010;
    cos[158] = 32'b1111111111111111_0001001010100101;
    cos[159] = 32'b1111111111111111_0001000100000001;
    cos[160] = 32'b1111111111111111_0000111101110001;
    cos[161] = 32'b1111111111111111_0000110111110011;
    cos[162] = 32'b1111111111111111_0000110010001000;
    cos[163] = 32'b1111111111111111_0000101100110000;
    cos[164] = 32'b1111111111111111_0000100111101011;
    cos[165] = 32'b1111111111111111_0000100010111010;
    cos[166] = 32'b1111111111111111_0000011110011011;
    cos[167] = 32'b1111111111111111_0000011010010000;
    cos[168] = 32'b1111111111111111_0000010110011001;
    cos[169] = 32'b1111111111111111_0000010010110101;
    cos[170] = 32'b1111111111111111_0000001111100100;
    cos[171] = 32'b1111111111111111_0000001100100111;
    cos[172] = 32'b1111111111111111_0000001001111110;
    cos[173] = 32'b1111111111111111_0000000111101001;
    cos[174] = 32'b1111111111111111_0000000101101000;
    cos[175] = 32'b1111111111111111_0000000011111010;
    cos[176] = 32'b1111111111111111_0000000010100000;
    cos[177] = 32'b1111111111111111_0000000001011010;
    cos[178] = 32'b1111111111111111_0000000000101000;
    cos[179] = 32'b1111111111111111_0000000000001010;
    cos[180] = 32'b1111111111111111_0000000000000000;


    PointsDrawLine[ 0][0] = 0; PointsDrawLine[ 0][1] = 1; 
    PointsDrawLine[ 1][0] = 1; PointsDrawLine[ 1][1] = 2; 
    PointsDrawLine[ 2][0] = 2; PointsDrawLine[ 2][1] = 3; 
    PointsDrawLine[ 3][0] = 3; PointsDrawLine[ 3][1] = 0; 
    PointsDrawLine[ 4][0] = 4; PointsDrawLine[ 4][1] = 5; 
    PointsDrawLine[ 5][0] = 5; PointsDrawLine[ 5][1] = 6; 
    PointsDrawLine[ 6][0] = 6; PointsDrawLine[ 6][1] = 7; 
    PointsDrawLine[ 7][0] = 7; PointsDrawLine[ 7][1] = 4; 
    PointsDrawLine[ 8][0] = 0; PointsDrawLine[ 8][1] = 4;         
    PointsDrawLine[ 9][0] = 1; PointsDrawLine[ 9][1] = 5; 
    PointsDrawLine[10][0] = 2; PointsDrawLine[10][1] = 6; 
    PointsDrawLine[11][0] = 3; PointsDrawLine[11][1] = 7; 


    //0 = x                      //1 = y                      //2 = z
    VertexBuffer[0][0] = -VERTEX_POINT;   VertexBuffer[0][1] = -VERTEX_POINT;   VertexBuffer[0][2] = -VERTEX_POINT;
    VertexBuffer[1][0] =  VERTEX_POINT;   VertexBuffer[1][1] = -VERTEX_POINT;   VertexBuffer[1][2] = -VERTEX_POINT;
    VertexBuffer[2][0] =  VERTEX_POINT;   VertexBuffer[2][1] =  VERTEX_POINT;   VertexBuffer[2][2] = -VERTEX_POINT;
    VertexBuffer[3][0] = -VERTEX_POINT;   VertexBuffer[3][1] =  VERTEX_POINT;   VertexBuffer[3][2] = -VERTEX_POINT;
    VertexBuffer[4][0] = -VERTEX_POINT;   VertexBuffer[4][1] = -VERTEX_POINT;   VertexBuffer[4][2] =  VERTEX_POINT;
    VertexBuffer[5][0] =  VERTEX_POINT;   VertexBuffer[5][1] = -VERTEX_POINT;   VertexBuffer[5][2] =  VERTEX_POINT;
    VertexBuffer[6][0] =  VERTEX_POINT;   VertexBuffer[6][1] =  VERTEX_POINT;   VertexBuffer[6][2] =  VERTEX_POINT;
    VertexBuffer[7][0] = -VERTEX_POINT;   VertexBuffer[7][1] =  VERTEX_POINT;   VertexBuffer[7][2] =  VERTEX_POINT;

    //    //rotating Z
    if (ROTATE_AXIS == ROTATE_Z) begin
      for (integer vertNum = 0; vertNum < 8; vertNum++) begin

        sinTheta = sin[THETA];
        cosTheta = cos[THETA]; 

        //Checked: works
        cordX = VertexBuffer[vertNum][0]; 
        cordY = VertexBuffer[vertNum][1];     

        //Checked: works
        XsinTheta = cordX * sinTheta;
        XcosTheta = cordX * cosTheta;
        YcosTheta = cordY * cosTheta;
        YsinTheta = cordY * sinTheta;

        //Checked: works
        newCordX = XcosTheta[47:16] - YsinTheta[47:16]; //might want to delete: [__]
        newCordY = YcosTheta[47:16] + XsinTheta[47:16]; 

        //round the numbers
        RotatedVertexBuffer[vertNum][0] = newCordX;
        RotatedVertexBuffer[vertNum][1] = newCordY;
        RotatedVertexBuffer[vertNum][2] = VertexBuffer[vertNum][2];

      end
    end

    //         //rotating Y
    if (ROTATE_AXIS == ROTATE_Y) begin
      for (integer vertNum = 0; vertNum < 8; vertNum++) begin

        sinTheta = sin[THETA];
        cosTheta = cos[THETA]; 

        //Checked: works
        cordZ = VertexBuffer[vertNum][2]; 
        cordX = VertexBuffer[vertNum][0];     

        //Checked: works
        ZsinTheta = cordZ * sinTheta;
        ZcosTheta = cordZ * cosTheta;
        XcosTheta = cordX * cosTheta;
        XsinTheta = cordX * sinTheta;

        //Checked: works
        newCordX = XcosTheta[47:16] + ZsinTheta[47:16]; 
        newCordZ = ZcosTheta[47:16] - XsinTheta[47:16]; //might want to delete: [__]

        //round the numbers
        RotatedVertexBuffer[vertNum][0] = newCordX;
        RotatedVertexBuffer[vertNum][1] = VertexBuffer[vertNum][1];
        RotatedVertexBuffer[vertNum][2] = newCordZ;

      end
    end



    //rotating X
    if (ROTATE_AXIS == ROTATE_X) begin
      for (integer vertNum = 0; vertNum < 8; vertNum++) begin

        sinTheta = sin[THETA];
        cosTheta = cos[THETA]; 

        //Checked: works
        cordZ = VertexBuffer[vertNum][2]; 
        cordY = VertexBuffer[vertNum][1];     

        //Checked: works
        ZsinTheta = cordZ * sinTheta;
        ZcosTheta = cordZ * cosTheta;
        YcosTheta = cordY * cosTheta;
        YsinTheta = cordY * sinTheta;

        //Checked: works
        newCordY = YcosTheta[47:16] - ZsinTheta[47:16]; 
        newCordZ = ZcosTheta[47:16] + YsinTheta[47:16]; //might want to delete: [__]

        //round the numbers
        RotatedVertexBuffer[vertNum][0] = VertexBuffer[vertNum][0];
        RotatedVertexBuffer[vertNum][1] = newCordY;
        RotatedVertexBuffer[vertNum][2] = newCordZ;

      end
    end

    //ROTATE ALL
    if (ROTATE_AXIS == ROTATE_ALL) begin
      for (integer vertNum = 0; vertNum < 8; vertNum++) begin

        sinTheta = sin[THETA];
        cosTheta = cos[THETA]; 

        //Checked: works
        cordX = VertexBuffer[vertNum][0]; 
        cordY = VertexBuffer[vertNum][1];
        cordZ = VertexBuffer[vertNum][2];     

        //Checked: works
        XcosTheta = cordX * cosTheta;
        XsinTheta = cordX * sinTheta;
        YcosTheta = cordY * cosTheta;
        YsinTheta = cordY * sinTheta;
        ZsinTheta = cordZ * sinTheta;
        ZcosTheta = cordZ * cosTheta;

        //Checked: works
        newCordX = XcosTheta[47:16] + ZsinTheta[47:16]; 
        newCordY = YcosTheta[47:16] - ZsinTheta[47:16]; 
        newCordZ = ZcosTheta[47:16] + YsinTheta[47:16]; 

        //round the numbers
        RotatedVertexBuffer[vertNum][0] = newCordX;
        RotatedVertexBuffer[vertNum][1] = newCordY;
        RotatedVertexBuffer[vertNum][2] = newCordZ;

      end
    end  







    for (integer x = 0; x <= SIZE; x++) begin
      for (integer y = 0; y <= SIZE; y++) begin
        FrameBuffer[x][y] = 1'b0;
      end
    end

    for (integer i = 0; i < 12; i++) begin

      x1 = RotatedVertexBuffer[PointsDrawLine[i][0]][0];
      x2 = RotatedVertexBuffer[PointsDrawLine[i][1]][0];
      y1 = RotatedVertexBuffer[PointsDrawLine[i][0]][1];
      y2 = RotatedVertexBuffer[PointsDrawLine[i][1]][1];
      z1 = RotatedVertexBuffer[PointsDrawLine[i][0]][2];
      z2 = RotatedVertexBuffer[PointsDrawLine[i][1]][2];

      FrameBuffer[x1 + (SIZE/2)][y1 + (SIZE/2)] = 1'b1;
      FrameBuffer[x2 + (SIZE/2)][y2 + (SIZE/2)] = 1'b1;

      //get abolsute values of differnce of x
      dx = x2 - x1;
      if (dx < 0) begin
        dxAbs = -1 * dx;
      end
      else begin
        dxAbs = dx;
      end


      //get abolsute values of differnce of y
      dy = y2 - y1;
      if (dy < 0) begin
        dyAbs = -1 * dy;
      end
      else begin
        dyAbs = dy;
      end

      //get abolsute values of differnce of z
      dz = z2 - z1;
      if (dz < 0) begin
        dzAbs = -1 * dz;
      end
      else begin
        dzAbs = dz;
      end


      // set 's to 1 or -1
      //x
      if (x2 > x1) begin
        xs = 1; 
      end else begin
        xs = -1;
      end
      //y
      if (y2 > y1) begin
        ys = 1; 
      end else begin
        ys = -1;
      end
      //z
      if (z2 > z1) begin
        zs = 1; 
      end else begin
        zs = -1;
      end


      if (dxAbs >= dyAbs && dxAbs >= dzAbs) begin
        p1 = 2 * dyAbs - dxAbs;
        p2 = 2 * dyAbs - dxAbs; 
        while (x1 != x2) begin

          x1 += xs;
          if (p1 >= 0) begin 
            y1 += ys; 
            p1 -= 2 * dxAbs; 
          end
          if (p2 >= 0)begin 
            z1 += zs; 
            p2 -= 2 * dxAbs; 
          end
          p1 += 2 * dyAbs; 
          p2 += 2 * dzAbs; 

          FrameBuffer[x1 + (SIZE/2)][y1 + (SIZE/2)] = 1'b1;
        end
      end

      if (dyAbs >= dxAbs && dyAbs >= dzAbs) begin
        p1 = 2 * dxAbs - dyAbs;
        p2 = 2 * dzAbs - dyAbs;
       while (y1 != y2) begin
          y1 += ys;
          if (p1 >= 0) begin 
            x1 += xs; 
            p1 -= 2 * dyAbs; 
          end
          if (p2 >= 0)begin 
            z1 += zs; 
            p2 -= 2 * dyAbs; 
          end
          p1 += 2 * dxAbs; 
          p2 += 2 * dzAbs; 

          FrameBuffer[x1 + (SIZE/2)][y1 + (SIZE/2)] = 1'b1;
        end
      end
      //z
      else begin
        p1 = 2 * dyAbs - dzAbs;
        p2 = 2 * dxAbs - dzAbs;
        while(z1 != z2) begin
          z1 += zs;
          if (p1 >= 0) begin 
            y1 += ys; 
            p1 -= 2 * dzAbs; 
          end
          if (p2 >= 0)begin 
            x1 += xs; 
            p2 -= 2 * dzAbs; 
          end
          p1 += 2 * dyAbs; 
          p2 += 2 * dxAbs; 

          FrameBuffer[x1 + (SIZE/2)][y1 + (SIZE/2)] = 1'b1;
        end
      end
    end
  end

endmodule
